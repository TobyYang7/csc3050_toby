// `include "alu.v"

`timescale 1ns/1ps

module test_alu();
    reg[31:0] instruction, regA, regB;
    wire[31:0] result;
    wire[2:0] flags;

    alu test(
        .instruction (instruction),
        .regA (regA),
        .regB (regB),
        .result (result), 
        .flags (flags)
    );

    initial begin
        $monitor("Time: %3d.\n Instruction: %32b\n regA: %32b, regB: %32b\n result: %32b, flags: %3b\n",
        $time, instruction, regA, regB, result, flags);

        // add
        #1
        $display("add");
        instruction = 32'b000000_00000_00001_00000_00000_100000; //000000 00000 00001 00000 00000 100000
        regA = 32'b000000_00000_00000_00000_00000_000001;
        regB = 32'b000000_00000_00000_00000_00000_000001; 

        // add with overflow-positive
        #1
        $display("add with overflow-positive");
        instruction = 32'b000000_00000_00001_00000_00000_100000;
        regA = 32'b01111111_11111111_11111111_11111111;
        regB = 32'b01111111_11111111_11111111_11111111;

        // add with overflow-negative
        #1
        $display("add with overflow-negative");
        instruction = 32'b000000_00000_00001_00000_00000_100000;
        regA = 32'b10000000_00000000_00000000_00000000;
        regB = 32'b10000000_00000000_00000000_00000000;

        // addi
        #1
        $display("addi");
        instruction = 32'b001000_00001_00000_01111_11111_111111;
        regA = 32'b01111111_11111111_11111111_11111111;
        regB = 32'b000000_00000_00000_00000_00000_000001;

        // addi with overflow
        #1
        $display("addi with overflow");
        instruction = 32'b001000_00000_00001_01111_11111_111111;
        regA = 32'b01111111_11111111_11111111_11111111;
        regB = 32'b000000_00000_00000_00000_00000_000001;

        // addu
        #1
        $display("addu");
        instruction = 32'b000000_00000_00001_00000_00000_100001;
        regA = 32'b1;
        regB = 32'b11111111_11111111_11111111_11111110;

        // addiu
        #1
        $display("addiu");
        instruction = 32'b001001_00000_00001_0111111111111111;
        regA = 32'b01111111_11111111_11111111_11111111;
        regB = 32'b1;

        // sub
        #1
        $display("sub");
        instruction = 32'b000000_00000_00001_00000_00000_100010;
        regA = 32'b1;
        regB = 32'b1;

        // sub with overflow-positive
        #1
        $display("sub with overflow-positive");
        instruction = 32'b000000_00000_00001_00000_00000_100010;
        regA = 32'b01111111_11111111_11111111_11111111;
        regB = 32'b10000000_00000000_00000000_00000000;

        // sub with overflow-negative
        #1
        $display("sub with overflow-negative");
        instruction = 32'b000000_00000_00001_00000_00000_100010;
        regA = 32'b10000000_00000000_00000000_00000000;
        regB = 32'b01111111_11111111_11111111_11111111;

        // subu
        #1
        $display("subu");
        instruction = 32'b000000_00000_00001_00000_00000_100011;
        regA = 32'b10000000_00000000_00000000_00000000;
        regB = 32'b01111111_11111111_11111111_11111111;

        // and
        #1
        $display("and");
        instruction = 32'b000000_00000_00001_00000_00000_100100;
        regA = 32'b01111111_11111111_11111111_11111111;
        regB = 32'b00000000_00000000_00000000_11111111;

        // andi
        #1
        $display("andi");
        instruction = 32'b001100_00000_00001_00000_00011_111111;
        regA = 32'b01111111_11111111_11111111_11111111;
        regB = 32'b00000000_00000000_00000000_00000000;

        // nor
        #1
        $display("nor");
        instruction = 32'b000000_00000_00001_00000_00000_100111;
        regA = 32'b01111111_11111111_11111111_11111111;
        regB = 32'b00000000_00000000_00000000_11111111;

        // or
        #1
        $display("or");
        instruction = 32'b000000_00000_00001_00000_00000_100101;
        regA = 32'b01111111_11111111_11111111_11111111;
        regB = 32'b00000000_00000000_00000000_11111111;

        // ori
        #1
        $display("ori");
        instruction = 32'b001101_00000_00001_00000_00011_111111;
        regA = 32'b01111111_11111111_11111111_11111111;
        regB = 32'b11111111_11111111_11111111_11111110;

        // xor
        #1
        $display("xor");
        instruction = 32'b000000_00000_00001_00000_00000_100110;
        regA = 32'b01111111_11111111_11111111_11111111;
        regB = 32'b00000000_00000000_00000000_11111111;

        // ori
        #1
        $display("ori");
        instruction = 32'b001110_00000_00001_00000_00011_111111;
        regA = 32'b01111111_11111111_11111111_11111111;
        regB = 32'b11111111_11111111_11111111_11111110;

        // beq on equal
        #1
        $display("beq on equal");
        instruction = 32'b000100_00000_00001_00000_00000_000000;
        regA = 32'b00000000_00000000_00000000_00000001;
        regB = 32'b00000000_00000000_00000000_00000001;

        // beq on not equal
        #1
        $display("beq on not equal");
        instruction = 32'b000100_00000_00001_00000_00000_000000;
        regA = 32'b00000000_00000000_00000000_00000001;
        regB = 32'b00000000_00000000_00000000_00000000;

        // bne on equal
        #1
        $display("bne on equal");
        instruction = 32'b000101_00000_00001_00000_00000_000000;
        regA = 32'b00000000_00000000_00000000_00000001;
        regB = 32'b00000000_00000000_00000000_00000001;

        // bne on not equal
        #1
        $display("bne on not equal");
        instruction = 32'b000101_00000_00001_00000_00000_000000;
        regA = 32'b00000000_00000000_00000000_00000001;
        regB = 32'b00000000_00000000_00000000_00000000;

        // slt on less
        #1
        $display("slt on less");
        instruction = 32'b000000_00000_00001_00000_00000_101010;
        regA = 32'b11111111_11111111_11111111_11111111;
        regB = 32'b00000000_00000000_00000000_00000001;

        // slt on greater
        #1
        $display("slt on greater");
        instruction = 32'b000000_00000_00001_00000_00000_101010;
        regA = 32'b00000000_00000000_00000000_00000001;
        regB = 32'b00000000_00000000_00000000_00000000;

        // slti on less
        #1
        $display("slti on less");
        instruction = 32'b001010_00000_00001_01111_11111_111111;
        regA = 32'b11111111_11111111_11111111_11111111;
        regB = 32'b11111111_11111111_11111111_11111111;

        // slti on greater
        #1
        $display("slti on greater");
        instruction = 32'b001010_00000_00001_11111_11111_111111;
        regA = 32'b01111111_11111111_11111111_11111111;
        regB = 32'b00000000_00000000_00000000_00000000;

        // sltiu on less
        #1
        $display("sltiu on less");
        instruction = 32'b001011_00000_00001_11111_11111_111111;
        regA = 32'b00000000_00000000_00000000_00000000;
        regB = 32'b00000000_00000000_00000000_00000001;

        // sltiu on greater
        #1
        $display("sltiu on greater");
        instruction = 32'b001011_00000_00001_11111_11111_111111;
        regA = 32'b11111111_11111111_11111111_11111111;
        regB = 32'b00000000_00000000_00000000_00000000;

        // sltu on less
        #1
        $display("sltu on less");
        instruction = 32'b000000_00000_00001_00000_00000_101011;
        regA = 32'b00000000_00000000_00000000_00000000;
        regB = 32'b00000000_00000000_00000000_00000001;

        // sltu on greater
        #1
        $display("sltu on greater");
        instruction = 32'b000000_00000_00001_00000_00000_101011;
        regA = 32'b11111111_11111111_11111111_11111111;
        regB = 32'b00000000_00000000_00000000_00000000;

        // lw
        #1
        $display("lw");
        instruction = 32'b100011_00000_00001_00000_00000_000000;
        regA = 32'b00000000_00000000_00000000_00000001;
        regB = 32'b00000000_00000000_00000000_00000000;

        // sw
        #1
        $display("sw");
        instruction = 32'b101011_00000_00001_00000_00000_000000;
        regA = 32'b00000000_00000000_00000000_00000001;
        regB = 32'b00000000_00000000_00000000_00000000;

        // sll
        #1
        $display("sll");
        instruction = 32'b000000_00000_00001_00000_00100_000000;
        regA = 32'b00000000_00000000_00000000_00000000;
        regB = 32'b11111111_11111111_11111111_11111111;

        // sllv
        #1
        $display("sllv");
        instruction = 32'b000000_00000_00001_00000_00100_000100;
        regA = 32'b00000000_00000000_00000000_00000100;
        regB = 32'b11111111_11111111_11111111_11111111;

        // srl
        #1
        $display("srl");
        instruction = 32'b000000_00000_00001_00000_00100_000010;
        regA = 32'b00000000_00000000_00000000_00000000;
        regB = 32'b11111111_11111111_11111111_11111111;

        // srlv
        #1
        $display("srlv");
        instruction = 32'b000000_00000_00001_00000_00100_000110;
        regA = 32'b00000000_00000000_00000000_00000100;
        regB = 32'b11111111_11111111_11111111_11111111;

        // sra
        #1
        $display("sra");
        instruction = 32'b000000_00000_00001_00000_00100_000011;
        regA = 32'b00000000_00000000_00000000_00000000;
        regB = 32'b10000000_11111111_11111111_11111111;

        // srav
        #1
        $display("srav");
        instruction = 32'b000000_00000_00001_00000_00100_000111;
        regA = 32'b00000000_00000000_00000000_00000100;
        regB = 32'b10000000_11111111_11111111_11111111;
    end

endmodule
